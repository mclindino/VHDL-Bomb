library verilog;
use verilog.vl_types.all;
entity Bombeador_vlg_vec_tst is
end Bombeador_vlg_vec_tst;
