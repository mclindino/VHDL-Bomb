library verilog;
use verilog.vl_types.all;
entity Bombeador_vlg_check_tst is
    port(
        clock_end       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Bombeador_vlg_check_tst;
